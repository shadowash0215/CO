module string_to_print #(parameter str_idx_end=1436) (
  input  [11:0] str_idx    ,
  output [ 7:0] data       ,
  input  [31:0] pc_if      ,
  input  [31:0] inst_if    ,
  input  [31:0] pc_id      ,
  input  [31:0] inst_id    ,
  input         valid_id   ,
  input  [31:0] x0         ,
  input  [31:0] ra         ,
  input  [31:0] sp         ,
  input  [31:0] gp         ,
  input  [31:0] tp         ,
  input  [31:0] t0         ,
  input  [31:0] t1         ,
  input  [31:0] t2         ,
  input  [31:0] s0         ,
  input  [31:0] s1         ,
  input  [31:0] a0         ,
  input  [31:0] a1         ,
  input  [31:0] a2         ,
  input  [31:0] a3         ,
  input  [31:0] a4         ,
  input  [31:0] a5         ,
  input  [31:0] a6         ,
  input  [31:0] a7         ,
  input  [31:0] s2         ,
  input  [31:0] s3         ,
  input  [31:0] s4         ,
  input  [31:0] s5         ,
  input  [31:0] s6         ,
  input  [31:0] s7         ,
  input  [31:0] s8         ,
  input  [31:0] s9         ,
  input  [31:0] s10        ,
  input  [31:0] s11        ,
  input  [31:0] t3         ,
  input  [31:0] t4         ,
  input  [31:0] t5         ,
  input  [31:0] t6         ,
  input  [31:0] pc_ex      ,
  input  [31:0] inst_ex    ,
  input         valid_ex   ,
  input  [ 4:0] rd_ex      ,
  input  [ 4:0] rs1        ,
  input  [ 4:0] rs2        ,
  input  [31:0] rs1_val    ,
  input  [31:0] rs2_val    ,
  input         reg_wen_ex ,
  input         is_imm     ,
  input  [31:0] imm        ,
  input         mem_wen_ex ,
  input         mem_ren_ex ,
  input         is_branch  ,
  input         is_jal_ex  ,
  input         is_jalr_ex ,
  input         is_auipc   ,
  input         is_lui     ,
  input  [ 3:0] alu_ctrl   ,
  input  [ 2:0] cmp_ctrl   ,
  input  [31:0] pc_mem     ,
  input  [31:0] inst_mem   ,
  input         valid_mem  ,
  input  [ 4:0] rd_mem     ,
  input         reg_wen_mem,
  input  [31:0] mem_w_data ,
  input  [31:0] alu_res    ,
  input         mem_wen_mem,
  input         mem_ren_mem,
  input         is_jal_mem ,
  input         is_jalr_mem,
  input  [31:0] pc_wb      ,
  input  [31:0] inst_wb    ,
  input         valid_wb   ,
  input  [ 4:0] rd_wb      ,
  input         reg_wen_wb ,
  input  [31:0] reg_w_data
);

  wire[7:0] str_print[str_idx_end-1:0];
  assign data = str_print[str_idx];

  // Value for constant part
  assign str_print[0]    = 8'h52;
  assign str_print[1]    = 8'h56;
  assign str_print[2]    = 8'h33;
  assign str_print[3]    = 8'h32;
  assign str_print[4]    = 8'h49;
  assign str_print[5]    = 8'h20;
  assign str_print[6]    = 8'h50;
  assign str_print[7]    = 8'h69;
  assign str_print[8]    = 8'h70;
  assign str_print[9]    = 8'h65;
  assign str_print[10]   = 8'h6C;
  assign str_print[11]   = 8'h69;
  assign str_print[12]   = 8'h6E;
  assign str_print[13]   = 8'h65;
  assign str_print[14]   = 8'h64;
  assign str_print[15]   = 8'h20;
  assign str_print[16]   = 8'h43;
  assign str_print[17]   = 8'h50;
  assign str_print[18]   = 8'h55;
  assign str_print[19]   = 8'h0A;
  assign str_print[20]   = 8'h0D;
  assign str_print[21]   = 8'h0A;
  assign str_print[22]   = 8'h0D;
  assign str_print[23]   = 8'h3D;
  assign str_print[24]   = 8'h3D;
  assign str_print[25]   = 8'h3D;
  assign str_print[26]   = 8'h3D;
  assign str_print[27]   = 8'h3D;
  assign str_print[28]   = 8'h3D;
  assign str_print[29]   = 8'h3D;
  assign str_print[30]   = 8'h3D;
  assign str_print[31]   = 8'h3D;
  assign str_print[32]   = 8'h3D;
  assign str_print[33]   = 8'h3D;
  assign str_print[34]   = 8'h3D;
  assign str_print[35]   = 8'h3D;
  assign str_print[36]   = 8'h3D;
  assign str_print[37]   = 8'h3D;
  assign str_print[38]   = 8'h3D;
  assign str_print[39]   = 8'h3D;
  assign str_print[40]   = 8'h3D;
  assign str_print[41]   = 8'h3D;
  assign str_print[42]   = 8'h3D;
  assign str_print[43]   = 8'h3D;
  assign str_print[44]   = 8'h3D;
  assign str_print[45]   = 8'h3D;
  assign str_print[46]   = 8'h3D;
  assign str_print[47]   = 8'h3D;
  assign str_print[48]   = 8'h3D;
  assign str_print[49]   = 8'h3D;
  assign str_print[50]   = 8'h3D;
  assign str_print[51]   = 8'h3D;
  assign str_print[52]   = 8'h3D;
  assign str_print[53]   = 8'h3D;
  assign str_print[54]   = 8'h3D;
  assign str_print[55]   = 8'h3D;
  assign str_print[56]   = 8'h3D;
  assign str_print[57]   = 8'h3D;
  assign str_print[58]   = 8'h3D;
  assign str_print[59]   = 8'h3D;
  assign str_print[60]   = 8'h3D;
  assign str_print[61]   = 8'h20;
  assign str_print[62]   = 8'h49;
  assign str_print[63]   = 8'h66;
  assign str_print[64]   = 8'h20;
  assign str_print[65]   = 8'h3D;
  assign str_print[66]   = 8'h3D;
  assign str_print[67]   = 8'h3D;
  assign str_print[68]   = 8'h3D;
  assign str_print[69]   = 8'h3D;
  assign str_print[70]   = 8'h3D;
  assign str_print[71]   = 8'h3D;
  assign str_print[72]   = 8'h3D;
  assign str_print[73]   = 8'h3D;
  assign str_print[74]   = 8'h3D;
  assign str_print[75]   = 8'h3D;
  assign str_print[76]   = 8'h3D;
  assign str_print[77]   = 8'h3D;
  assign str_print[78]   = 8'h3D;
  assign str_print[79]   = 8'h3D;
  assign str_print[80]   = 8'h3D;
  assign str_print[81]   = 8'h3D;
  assign str_print[82]   = 8'h3D;
  assign str_print[83]   = 8'h3D;
  assign str_print[84]   = 8'h3D;
  assign str_print[85]   = 8'h3D;
  assign str_print[86]   = 8'h3D;
  assign str_print[87]   = 8'h3D;
  assign str_print[88]   = 8'h3D;
  assign str_print[89]   = 8'h3D;
  assign str_print[90]   = 8'h3D;
  assign str_print[91]   = 8'h3D;
  assign str_print[92]   = 8'h3D;
  assign str_print[93]   = 8'h3D;
  assign str_print[94]   = 8'h3D;
  assign str_print[95]   = 8'h3D;
  assign str_print[96]   = 8'h3D;
  assign str_print[97]   = 8'h3D;
  assign str_print[98]   = 8'h3D;
  assign str_print[99]   = 8'h3D;
  assign str_print[100]  = 8'h3D;
  assign str_print[101]  = 8'h3D;
  assign str_print[102]  = 8'h3D;
  assign str_print[103]  = 8'h3D;
  assign str_print[104]  = 8'h0A;
  assign str_print[105]  = 8'h0D;
  assign str_print[106]  = 8'h70;
  assign str_print[107]  = 8'h63;
  assign str_print[108]  = 8'h3A;
  assign str_print[109]  = 8'h20;
  assign str_print[118]  = 8'h09;
  assign str_print[119]  = 8'h69;
  assign str_print[120]  = 8'h6E;
  assign str_print[121]  = 8'h73;
  assign str_print[122]  = 8'h74;
  assign str_print[123]  = 8'h3A;
  assign str_print[124]  = 8'h20;
  assign str_print[133]  = 8'h0A;
  assign str_print[134]  = 8'h0D;
  assign str_print[135]  = 8'h3D;
  assign str_print[136]  = 8'h3D;
  assign str_print[137]  = 8'h3D;
  assign str_print[138]  = 8'h3D;
  assign str_print[139]  = 8'h3D;
  assign str_print[140]  = 8'h3D;
  assign str_print[141]  = 8'h3D;
  assign str_print[142]  = 8'h3D;
  assign str_print[143]  = 8'h3D;
  assign str_print[144]  = 8'h3D;
  assign str_print[145]  = 8'h3D;
  assign str_print[146]  = 8'h3D;
  assign str_print[147]  = 8'h3D;
  assign str_print[148]  = 8'h3D;
  assign str_print[149]  = 8'h3D;
  assign str_print[150]  = 8'h3D;
  assign str_print[151]  = 8'h3D;
  assign str_print[152]  = 8'h3D;
  assign str_print[153]  = 8'h3D;
  assign str_print[154]  = 8'h3D;
  assign str_print[155]  = 8'h3D;
  assign str_print[156]  = 8'h3D;
  assign str_print[157]  = 8'h3D;
  assign str_print[158]  = 8'h3D;
  assign str_print[159]  = 8'h3D;
  assign str_print[160]  = 8'h3D;
  assign str_print[161]  = 8'h3D;
  assign str_print[162]  = 8'h3D;
  assign str_print[163]  = 8'h3D;
  assign str_print[164]  = 8'h3D;
  assign str_print[165]  = 8'h3D;
  assign str_print[166]  = 8'h3D;
  assign str_print[167]  = 8'h3D;
  assign str_print[168]  = 8'h3D;
  assign str_print[169]  = 8'h3D;
  assign str_print[170]  = 8'h3D;
  assign str_print[171]  = 8'h3D;
  assign str_print[172]  = 8'h3D;
  assign str_print[173]  = 8'h20;
  assign str_print[174]  = 8'h49;
  assign str_print[175]  = 8'h64;
  assign str_print[176]  = 8'h20;
  assign str_print[177]  = 8'h3D;
  assign str_print[178]  = 8'h3D;
  assign str_print[179]  = 8'h3D;
  assign str_print[180]  = 8'h3D;
  assign str_print[181]  = 8'h3D;
  assign str_print[182]  = 8'h3D;
  assign str_print[183]  = 8'h3D;
  assign str_print[184]  = 8'h3D;
  assign str_print[185]  = 8'h3D;
  assign str_print[186]  = 8'h3D;
  assign str_print[187]  = 8'h3D;
  assign str_print[188]  = 8'h3D;
  assign str_print[189]  = 8'h3D;
  assign str_print[190]  = 8'h3D;
  assign str_print[191]  = 8'h3D;
  assign str_print[192]  = 8'h3D;
  assign str_print[193]  = 8'h3D;
  assign str_print[194]  = 8'h3D;
  assign str_print[195]  = 8'h3D;
  assign str_print[196]  = 8'h3D;
  assign str_print[197]  = 8'h3D;
  assign str_print[198]  = 8'h3D;
  assign str_print[199]  = 8'h3D;
  assign str_print[200]  = 8'h3D;
  assign str_print[201]  = 8'h3D;
  assign str_print[202]  = 8'h3D;
  assign str_print[203]  = 8'h3D;
  assign str_print[204]  = 8'h3D;
  assign str_print[205]  = 8'h3D;
  assign str_print[206]  = 8'h3D;
  assign str_print[207]  = 8'h3D;
  assign str_print[208]  = 8'h3D;
  assign str_print[209]  = 8'h3D;
  assign str_print[210]  = 8'h3D;
  assign str_print[211]  = 8'h3D;
  assign str_print[212]  = 8'h3D;
  assign str_print[213]  = 8'h3D;
  assign str_print[214]  = 8'h3D;
  assign str_print[215]  = 8'h3D;
  assign str_print[216]  = 8'h0A;
  assign str_print[217]  = 8'h0D;
  assign str_print[218]  = 8'h70;
  assign str_print[219]  = 8'h63;
  assign str_print[220]  = 8'h3A;
  assign str_print[221]  = 8'h20;
  assign str_print[230]  = 8'h09;
  assign str_print[231]  = 8'h69;
  assign str_print[232]  = 8'h6E;
  assign str_print[233]  = 8'h73;
  assign str_print[234]  = 8'h74;
  assign str_print[235]  = 8'h3A;
  assign str_print[236]  = 8'h20;
  assign str_print[245]  = 8'h09;
  assign str_print[246]  = 8'h76;
  assign str_print[247]  = 8'h61;
  assign str_print[248]  = 8'h6C;
  assign str_print[249]  = 8'h69;
  assign str_print[250]  = 8'h64;
  assign str_print[251]  = 8'h3A;
  assign str_print[252]  = 8'h20;
  assign str_print[254]  = 8'h0A;
  assign str_print[255]  = 8'h0D;
  assign str_print[256]  = 8'h78;
  assign str_print[257]  = 8'h30;
  assign str_print[258]  = 8'h3A;
  assign str_print[259]  = 8'h20;
  assign str_print[268]  = 8'h09;
  assign str_print[269]  = 8'h72;
  assign str_print[270]  = 8'h61;
  assign str_print[271]  = 8'h3A;
  assign str_print[272]  = 8'h20;
  assign str_print[281]  = 8'h09;
  assign str_print[282]  = 8'h73;
  assign str_print[283]  = 8'h70;
  assign str_print[284]  = 8'h3A;
  assign str_print[285]  = 8'h20;
  assign str_print[294]  = 8'h09;
  assign str_print[295]  = 8'h67;
  assign str_print[296]  = 8'h70;
  assign str_print[297]  = 8'h3A;
  assign str_print[298]  = 8'h20;
  assign str_print[307]  = 8'h09;
  assign str_print[308]  = 8'h74;
  assign str_print[309]  = 8'h70;
  assign str_print[310]  = 8'h3A;
  assign str_print[311]  = 8'h20;
  assign str_print[320]  = 8'h0A;
  assign str_print[321]  = 8'h0D;
  assign str_print[322]  = 8'h74;
  assign str_print[323]  = 8'h30;
  assign str_print[324]  = 8'h3A;
  assign str_print[325]  = 8'h20;
  assign str_print[334]  = 8'h09;
  assign str_print[335]  = 8'h74;
  assign str_print[336]  = 8'h31;
  assign str_print[337]  = 8'h3A;
  assign str_print[338]  = 8'h20;
  assign str_print[347]  = 8'h09;
  assign str_print[348]  = 8'h74;
  assign str_print[349]  = 8'h32;
  assign str_print[350]  = 8'h3A;
  assign str_print[351]  = 8'h20;
  assign str_print[360]  = 8'h09;
  assign str_print[361]  = 8'h73;
  assign str_print[362]  = 8'h30;
  assign str_print[363]  = 8'h3A;
  assign str_print[364]  = 8'h20;
  assign str_print[373]  = 8'h09;
  assign str_print[374]  = 8'h73;
  assign str_print[375]  = 8'h31;
  assign str_print[376]  = 8'h3A;
  assign str_print[377]  = 8'h20;
  assign str_print[386]  = 8'h0A;
  assign str_print[387]  = 8'h0D;
  assign str_print[388]  = 8'h61;
  assign str_print[389]  = 8'h30;
  assign str_print[390]  = 8'h3A;
  assign str_print[391]  = 8'h20;
  assign str_print[400]  = 8'h09;
  assign str_print[401]  = 8'h61;
  assign str_print[402]  = 8'h31;
  assign str_print[403]  = 8'h3A;
  assign str_print[404]  = 8'h20;
  assign str_print[413]  = 8'h09;
  assign str_print[414]  = 8'h61;
  assign str_print[415]  = 8'h32;
  assign str_print[416]  = 8'h3A;
  assign str_print[417]  = 8'h20;
  assign str_print[426]  = 8'h09;
  assign str_print[427]  = 8'h61;
  assign str_print[428]  = 8'h33;
  assign str_print[429]  = 8'h3A;
  assign str_print[430]  = 8'h20;
  assign str_print[439]  = 8'h09;
  assign str_print[440]  = 8'h61;
  assign str_print[441]  = 8'h34;
  assign str_print[442]  = 8'h3A;
  assign str_print[443]  = 8'h20;
  assign str_print[452]  = 8'h0A;
  assign str_print[453]  = 8'h0D;
  assign str_print[454]  = 8'h61;
  assign str_print[455]  = 8'h35;
  assign str_print[456]  = 8'h3A;
  assign str_print[457]  = 8'h20;
  assign str_print[466]  = 8'h09;
  assign str_print[467]  = 8'h61;
  assign str_print[468]  = 8'h36;
  assign str_print[469]  = 8'h3A;
  assign str_print[470]  = 8'h20;
  assign str_print[479]  = 8'h09;
  assign str_print[480]  = 8'h61;
  assign str_print[481]  = 8'h37;
  assign str_print[482]  = 8'h3A;
  assign str_print[483]  = 8'h20;
  assign str_print[492]  = 8'h09;
  assign str_print[493]  = 8'h73;
  assign str_print[494]  = 8'h32;
  assign str_print[495]  = 8'h3A;
  assign str_print[496]  = 8'h20;
  assign str_print[505]  = 8'h09;
  assign str_print[506]  = 8'h73;
  assign str_print[507]  = 8'h33;
  assign str_print[508]  = 8'h3A;
  assign str_print[509]  = 8'h20;
  assign str_print[518]  = 8'h0A;
  assign str_print[519]  = 8'h0D;
  assign str_print[520]  = 8'h73;
  assign str_print[521]  = 8'h34;
  assign str_print[522]  = 8'h3A;
  assign str_print[523]  = 8'h20;
  assign str_print[532]  = 8'h09;
  assign str_print[533]  = 8'h73;
  assign str_print[534]  = 8'h35;
  assign str_print[535]  = 8'h3A;
  assign str_print[536]  = 8'h20;
  assign str_print[545]  = 8'h09;
  assign str_print[546]  = 8'h73;
  assign str_print[547]  = 8'h36;
  assign str_print[548]  = 8'h3A;
  assign str_print[549]  = 8'h20;
  assign str_print[558]  = 8'h09;
  assign str_print[559]  = 8'h73;
  assign str_print[560]  = 8'h37;
  assign str_print[561]  = 8'h3A;
  assign str_print[562]  = 8'h20;
  assign str_print[571]  = 8'h09;
  assign str_print[572]  = 8'h73;
  assign str_print[573]  = 8'h38;
  assign str_print[574]  = 8'h3A;
  assign str_print[575]  = 8'h20;
  assign str_print[584]  = 8'h0A;
  assign str_print[585]  = 8'h0D;
  assign str_print[586]  = 8'h73;
  assign str_print[587]  = 8'h39;
  assign str_print[588]  = 8'h3A;
  assign str_print[589]  = 8'h20;
  assign str_print[598]  = 8'h09;
  assign str_print[599]  = 8'h73;
  assign str_print[600]  = 8'h31;
  assign str_print[601]  = 8'h30;
  assign str_print[602]  = 8'h3A;
  assign str_print[611]  = 8'h09;
  assign str_print[612]  = 8'h73;
  assign str_print[613]  = 8'h31;
  assign str_print[614]  = 8'h31;
  assign str_print[615]  = 8'h3A;
  assign str_print[624]  = 8'h09;
  assign str_print[625]  = 8'h74;
  assign str_print[626]  = 8'h33;
  assign str_print[627]  = 8'h3A;
  assign str_print[628]  = 8'h20;
  assign str_print[637]  = 8'h09;
  assign str_print[638]  = 8'h74;
  assign str_print[639]  = 8'h34;
  assign str_print[640]  = 8'h3A;
  assign str_print[641]  = 8'h20;
  assign str_print[650]  = 8'h0A;
  assign str_print[651]  = 8'h0D;
  assign str_print[652]  = 8'h74;
  assign str_print[653]  = 8'h35;
  assign str_print[654]  = 8'h3A;
  assign str_print[655]  = 8'h20;
  assign str_print[664]  = 8'h09;
  assign str_print[665]  = 8'h74;
  assign str_print[666]  = 8'h36;
  assign str_print[667]  = 8'h3A;
  assign str_print[668]  = 8'h20;
  assign str_print[677]  = 8'h0A;
  assign str_print[678]  = 8'h0D;
  assign str_print[679]  = 8'h3D;
  assign str_print[680]  = 8'h3D;
  assign str_print[681]  = 8'h3D;
  assign str_print[682]  = 8'h3D;
  assign str_print[683]  = 8'h3D;
  assign str_print[684]  = 8'h3D;
  assign str_print[685]  = 8'h3D;
  assign str_print[686]  = 8'h3D;
  assign str_print[687]  = 8'h3D;
  assign str_print[688]  = 8'h3D;
  assign str_print[689]  = 8'h3D;
  assign str_print[690]  = 8'h3D;
  assign str_print[691]  = 8'h3D;
  assign str_print[692]  = 8'h3D;
  assign str_print[693]  = 8'h3D;
  assign str_print[694]  = 8'h3D;
  assign str_print[695]  = 8'h3D;
  assign str_print[696]  = 8'h3D;
  assign str_print[697]  = 8'h3D;
  assign str_print[698]  = 8'h3D;
  assign str_print[699]  = 8'h3D;
  assign str_print[700]  = 8'h3D;
  assign str_print[701]  = 8'h3D;
  assign str_print[702]  = 8'h3D;
  assign str_print[703]  = 8'h3D;
  assign str_print[704]  = 8'h3D;
  assign str_print[705]  = 8'h3D;
  assign str_print[706]  = 8'h3D;
  assign str_print[707]  = 8'h3D;
  assign str_print[708]  = 8'h3D;
  assign str_print[709]  = 8'h3D;
  assign str_print[710]  = 8'h3D;
  assign str_print[711]  = 8'h3D;
  assign str_print[712]  = 8'h3D;
  assign str_print[713]  = 8'h3D;
  assign str_print[714]  = 8'h3D;
  assign str_print[715]  = 8'h3D;
  assign str_print[716]  = 8'h3D;
  assign str_print[717]  = 8'h20;
  assign str_print[718]  = 8'h45;
  assign str_print[719]  = 8'h78;
  assign str_print[720]  = 8'h20;
  assign str_print[721]  = 8'h3D;
  assign str_print[722]  = 8'h3D;
  assign str_print[723]  = 8'h3D;
  assign str_print[724]  = 8'h3D;
  assign str_print[725]  = 8'h3D;
  assign str_print[726]  = 8'h3D;
  assign str_print[727]  = 8'h3D;
  assign str_print[728]  = 8'h3D;
  assign str_print[729]  = 8'h3D;
  assign str_print[730]  = 8'h3D;
  assign str_print[731]  = 8'h3D;
  assign str_print[732]  = 8'h3D;
  assign str_print[733]  = 8'h3D;
  assign str_print[734]  = 8'h3D;
  assign str_print[735]  = 8'h3D;
  assign str_print[736]  = 8'h3D;
  assign str_print[737]  = 8'h3D;
  assign str_print[738]  = 8'h3D;
  assign str_print[739]  = 8'h3D;
  assign str_print[740]  = 8'h3D;
  assign str_print[741]  = 8'h3D;
  assign str_print[742]  = 8'h3D;
  assign str_print[743]  = 8'h3D;
  assign str_print[744]  = 8'h3D;
  assign str_print[745]  = 8'h3D;
  assign str_print[746]  = 8'h3D;
  assign str_print[747]  = 8'h3D;
  assign str_print[748]  = 8'h3D;
  assign str_print[749]  = 8'h3D;
  assign str_print[750]  = 8'h3D;
  assign str_print[751]  = 8'h3D;
  assign str_print[752]  = 8'h3D;
  assign str_print[753]  = 8'h3D;
  assign str_print[754]  = 8'h3D;
  assign str_print[755]  = 8'h3D;
  assign str_print[756]  = 8'h3D;
  assign str_print[757]  = 8'h3D;
  assign str_print[758]  = 8'h3D;
  assign str_print[759]  = 8'h3D;
  assign str_print[760]  = 8'h0A;
  assign str_print[761]  = 8'h0D;
  assign str_print[762]  = 8'h70;
  assign str_print[763]  = 8'h63;
  assign str_print[764]  = 8'h3A;
  assign str_print[765]  = 8'h20;
  assign str_print[774]  = 8'h09;
  assign str_print[775]  = 8'h69;
  assign str_print[776]  = 8'h6E;
  assign str_print[777]  = 8'h73;
  assign str_print[778]  = 8'h74;
  assign str_print[779]  = 8'h3A;
  assign str_print[780]  = 8'h20;
  assign str_print[789]  = 8'h09;
  assign str_print[790]  = 8'h76;
  assign str_print[791]  = 8'h61;
  assign str_print[792]  = 8'h6C;
  assign str_print[793]  = 8'h69;
  assign str_print[794]  = 8'h64;
  assign str_print[795]  = 8'h3A;
  assign str_print[796]  = 8'h20;
  assign str_print[798]  = 8'h0A;
  assign str_print[799]  = 8'h0D;
  assign str_print[800]  = 8'h72;
  assign str_print[801]  = 8'h64;
  assign str_print[802]  = 8'h3A;
  assign str_print[803]  = 8'h20;
  assign str_print[804]  = 8'h20;
  assign str_print[807]  = 8'h09;
  assign str_print[808]  = 8'h72;
  assign str_print[809]  = 8'h73;
  assign str_print[810]  = 8'h31;
  assign str_print[811]  = 8'h3A;
  assign str_print[812]  = 8'h20;
  assign str_print[815]  = 8'h09;
  assign str_print[816]  = 8'h72;
  assign str_print[817]  = 8'h73;
  assign str_print[818]  = 8'h32;
  assign str_print[819]  = 8'h3A;
  assign str_print[820]  = 8'h20;
  assign str_print[823]  = 8'h09;
  assign str_print[824]  = 8'h72;
  assign str_print[825]  = 8'h73;
  assign str_print[826]  = 8'h31;
  assign str_print[827]  = 8'h5F;
  assign str_print[828]  = 8'h76;
  assign str_print[829]  = 8'h61;
  assign str_print[830]  = 8'h6C;
  assign str_print[831]  = 8'h3A;
  assign str_print[832]  = 8'h20;
  assign str_print[841]  = 8'h09;
  assign str_print[842]  = 8'h72;
  assign str_print[843]  = 8'h73;
  assign str_print[844]  = 8'h32;
  assign str_print[845]  = 8'h5F;
  assign str_print[846]  = 8'h76;
  assign str_print[847]  = 8'h61;
  assign str_print[848]  = 8'h6C;
  assign str_print[849]  = 8'h3A;
  assign str_print[850]  = 8'h20;
  assign str_print[859]  = 8'h09;
  assign str_print[860]  = 8'h72;
  assign str_print[861]  = 8'h65;
  assign str_print[862]  = 8'h67;
  assign str_print[863]  = 8'h5F;
  assign str_print[864]  = 8'h77;
  assign str_print[865]  = 8'h65;
  assign str_print[866]  = 8'h6E;
  assign str_print[867]  = 8'h3A;
  assign str_print[868]  = 8'h20;
  assign str_print[870]  = 8'h0A;
  assign str_print[871]  = 8'h0D;
  assign str_print[872]  = 8'h69;
  assign str_print[873]  = 8'h73;
  assign str_print[874]  = 8'h5F;
  assign str_print[875]  = 8'h69;
  assign str_print[876]  = 8'h6D;
  assign str_print[877]  = 8'h6D;
  assign str_print[878]  = 8'h3A;
  assign str_print[879]  = 8'h20;
  assign str_print[881]  = 8'h09;
  assign str_print[882]  = 8'h69;
  assign str_print[883]  = 8'h6D;
  assign str_print[884]  = 8'h6D;
  assign str_print[885]  = 8'h3A;
  assign str_print[886]  = 8'h20;
  assign str_print[895]  = 8'h0A;
  assign str_print[896]  = 8'h0D;
  assign str_print[897]  = 8'h6D;
  assign str_print[898]  = 8'h65;
  assign str_print[899]  = 8'h6D;
  assign str_print[900]  = 8'h5F;
  assign str_print[901]  = 8'h77;
  assign str_print[902]  = 8'h65;
  assign str_print[903]  = 8'h6E;
  assign str_print[904]  = 8'h3A;
  assign str_print[905]  = 8'h20;
  assign str_print[907]  = 8'h09;
  assign str_print[908]  = 8'h6D;
  assign str_print[909]  = 8'h65;
  assign str_print[910]  = 8'h6D;
  assign str_print[911]  = 8'h5F;
  assign str_print[912]  = 8'h72;
  assign str_print[913]  = 8'h65;
  assign str_print[914]  = 8'h6E;
  assign str_print[915]  = 8'h3A;
  assign str_print[916]  = 8'h20;
  assign str_print[918]  = 8'h09;
  assign str_print[919]  = 8'h69;
  assign str_print[920]  = 8'h73;
  assign str_print[921]  = 8'h5F;
  assign str_print[922]  = 8'h62;
  assign str_print[923]  = 8'h72;
  assign str_print[924]  = 8'h61;
  assign str_print[925]  = 8'h6E;
  assign str_print[926]  = 8'h63;
  assign str_print[927]  = 8'h68;
  assign str_print[928]  = 8'h3A;
  assign str_print[929]  = 8'h20;
  assign str_print[931]  = 8'h09;
  assign str_print[932]  = 8'h69;
  assign str_print[933]  = 8'h73;
  assign str_print[934]  = 8'h5F;
  assign str_print[935]  = 8'h6A;
  assign str_print[936]  = 8'h61;
  assign str_print[937]  = 8'h6C;
  assign str_print[938]  = 8'h3A;
  assign str_print[939]  = 8'h20;
  assign str_print[941]  = 8'h09;
  assign str_print[942]  = 8'h69;
  assign str_print[943]  = 8'h73;
  assign str_print[944]  = 8'h5F;
  assign str_print[945]  = 8'h6A;
  assign str_print[946]  = 8'h61;
  assign str_print[947]  = 8'h6C;
  assign str_print[948]  = 8'h72;
  assign str_print[949]  = 8'h3A;
  assign str_print[950]  = 8'h20;
  assign str_print[952]  = 8'h0A;
  assign str_print[953]  = 8'h0D;
  assign str_print[954]  = 8'h69;
  assign str_print[955]  = 8'h73;
  assign str_print[956]  = 8'h5F;
  assign str_print[957]  = 8'h61;
  assign str_print[958]  = 8'h75;
  assign str_print[959]  = 8'h69;
  assign str_print[960]  = 8'h70;
  assign str_print[961]  = 8'h63;
  assign str_print[962]  = 8'h3A;
  assign str_print[963]  = 8'h20;
  assign str_print[965]  = 8'h09;
  assign str_print[966]  = 8'h69;
  assign str_print[967]  = 8'h73;
  assign str_print[968]  = 8'h5F;
  assign str_print[969]  = 8'h6C;
  assign str_print[970]  = 8'h75;
  assign str_print[971]  = 8'h69;
  assign str_print[972]  = 8'h3A;
  assign str_print[973]  = 8'h20;
  assign str_print[975]  = 8'h09;
  assign str_print[976]  = 8'h61;
  assign str_print[977]  = 8'h6C;
  assign str_print[978]  = 8'h75;
  assign str_print[979]  = 8'h5F;
  assign str_print[980]  = 8'h63;
  assign str_print[981]  = 8'h74;
  assign str_print[982]  = 8'h72;
  assign str_print[983]  = 8'h6C;
  assign str_print[984]  = 8'h3A;
  assign str_print[985]  = 8'h20;
  assign str_print[987]  = 8'h09;
  assign str_print[988]  = 8'h63;
  assign str_print[989]  = 8'h6D;
  assign str_print[990]  = 8'h70;
  assign str_print[991]  = 8'h5F;
  assign str_print[992]  = 8'h63;
  assign str_print[993]  = 8'h74;
  assign str_print[994]  = 8'h72;
  assign str_print[995]  = 8'h6C;
  assign str_print[996]  = 8'h3A;
  assign str_print[997]  = 8'h20;
  assign str_print[999]  = 8'h0A;
  assign str_print[1000] = 8'h0D;
  assign str_print[1001] = 8'h3D;
  assign str_print[1002] = 8'h3D;
  assign str_print[1003] = 8'h3D;
  assign str_print[1004] = 8'h3D;
  assign str_print[1005] = 8'h3D;
  assign str_print[1006] = 8'h3D;
  assign str_print[1007] = 8'h3D;
  assign str_print[1008] = 8'h3D;
  assign str_print[1009] = 8'h3D;
  assign str_print[1010] = 8'h3D;
  assign str_print[1011] = 8'h3D;
  assign str_print[1012] = 8'h3D;
  assign str_print[1013] = 8'h3D;
  assign str_print[1014] = 8'h3D;
  assign str_print[1015] = 8'h3D;
  assign str_print[1016] = 8'h3D;
  assign str_print[1017] = 8'h3D;
  assign str_print[1018] = 8'h3D;
  assign str_print[1019] = 8'h3D;
  assign str_print[1020] = 8'h3D;
  assign str_print[1021] = 8'h3D;
  assign str_print[1022] = 8'h3D;
  assign str_print[1023] = 8'h3D;
  assign str_print[1024] = 8'h3D;
  assign str_print[1025] = 8'h3D;
  assign str_print[1026] = 8'h3D;
  assign str_print[1027] = 8'h3D;
  assign str_print[1028] = 8'h3D;
  assign str_print[1029] = 8'h3D;
  assign str_print[1030] = 8'h3D;
  assign str_print[1031] = 8'h3D;
  assign str_print[1032] = 8'h3D;
  assign str_print[1033] = 8'h3D;
  assign str_print[1034] = 8'h3D;
  assign str_print[1035] = 8'h3D;
  assign str_print[1036] = 8'h3D;
  assign str_print[1037] = 8'h3D;
  assign str_print[1038] = 8'h3D;
  assign str_print[1039] = 8'h20;
  assign str_print[1040] = 8'h4D;
  assign str_print[1041] = 8'h61;
  assign str_print[1042] = 8'h20;
  assign str_print[1043] = 8'h3D;
  assign str_print[1044] = 8'h3D;
  assign str_print[1045] = 8'h3D;
  assign str_print[1046] = 8'h3D;
  assign str_print[1047] = 8'h3D;
  assign str_print[1048] = 8'h3D;
  assign str_print[1049] = 8'h3D;
  assign str_print[1050] = 8'h3D;
  assign str_print[1051] = 8'h3D;
  assign str_print[1052] = 8'h3D;
  assign str_print[1053] = 8'h3D;
  assign str_print[1054] = 8'h3D;
  assign str_print[1055] = 8'h3D;
  assign str_print[1056] = 8'h3D;
  assign str_print[1057] = 8'h3D;
  assign str_print[1058] = 8'h3D;
  assign str_print[1059] = 8'h3D;
  assign str_print[1060] = 8'h3D;
  assign str_print[1061] = 8'h3D;
  assign str_print[1062] = 8'h3D;
  assign str_print[1063] = 8'h3D;
  assign str_print[1064] = 8'h3D;
  assign str_print[1065] = 8'h3D;
  assign str_print[1066] = 8'h3D;
  assign str_print[1067] = 8'h3D;
  assign str_print[1068] = 8'h3D;
  assign str_print[1069] = 8'h3D;
  assign str_print[1070] = 8'h3D;
  assign str_print[1071] = 8'h3D;
  assign str_print[1072] = 8'h3D;
  assign str_print[1073] = 8'h3D;
  assign str_print[1074] = 8'h3D;
  assign str_print[1075] = 8'h3D;
  assign str_print[1076] = 8'h3D;
  assign str_print[1077] = 8'h3D;
  assign str_print[1078] = 8'h3D;
  assign str_print[1079] = 8'h3D;
  assign str_print[1080] = 8'h3D;
  assign str_print[1081] = 8'h3D;
  assign str_print[1082] = 8'h0A;
  assign str_print[1083] = 8'h0D;
  assign str_print[1084] = 8'h70;
  assign str_print[1085] = 8'h63;
  assign str_print[1086] = 8'h3A;
  assign str_print[1087] = 8'h20;
  assign str_print[1096] = 8'h09;
  assign str_print[1097] = 8'h69;
  assign str_print[1098] = 8'h6E;
  assign str_print[1099] = 8'h73;
  assign str_print[1100] = 8'h74;
  assign str_print[1101] = 8'h3A;
  assign str_print[1102] = 8'h20;
  assign str_print[1111] = 8'h09;
  assign str_print[1112] = 8'h76;
  assign str_print[1113] = 8'h61;
  assign str_print[1114] = 8'h6C;
  assign str_print[1115] = 8'h69;
  assign str_print[1116] = 8'h64;
  assign str_print[1117] = 8'h3A;
  assign str_print[1118] = 8'h20;
  assign str_print[1120] = 8'h0A;
  assign str_print[1121] = 8'h0D;
  assign str_print[1122] = 8'h72;
  assign str_print[1123] = 8'h64;
  assign str_print[1124] = 8'h3A;
  assign str_print[1125] = 8'h20;
  assign str_print[1126] = 8'h20;
  assign str_print[1129] = 8'h09;
  assign str_print[1130] = 8'h72;
  assign str_print[1131] = 8'h65;
  assign str_print[1132] = 8'h67;
  assign str_print[1133] = 8'h5F;
  assign str_print[1134] = 8'h77;
  assign str_print[1135] = 8'h65;
  assign str_print[1136] = 8'h6E;
  assign str_print[1137] = 8'h3A;
  assign str_print[1138] = 8'h20;
  assign str_print[1140] = 8'h09;
  assign str_print[1141] = 8'h6D;
  assign str_print[1142] = 8'h65;
  assign str_print[1143] = 8'h6D;
  assign str_print[1144] = 8'h5F;
  assign str_print[1145] = 8'h77;
  assign str_print[1146] = 8'h5F;
  assign str_print[1147] = 8'h64;
  assign str_print[1148] = 8'h61;
  assign str_print[1149] = 8'h74;
  assign str_print[1150] = 8'h61;
  assign str_print[1151] = 8'h3A;
  assign str_print[1152] = 8'h20;
  assign str_print[1161] = 8'h09;
  assign str_print[1162] = 8'h61;
  assign str_print[1163] = 8'h6C;
  assign str_print[1164] = 8'h75;
  assign str_print[1165] = 8'h5F;
  assign str_print[1166] = 8'h72;
  assign str_print[1167] = 8'h65;
  assign str_print[1168] = 8'h73;
  assign str_print[1169] = 8'h3A;
  assign str_print[1170] = 8'h20;
  assign str_print[1179] = 8'h0A;
  assign str_print[1180] = 8'h0D;
  assign str_print[1181] = 8'h6D;
  assign str_print[1182] = 8'h65;
  assign str_print[1183] = 8'h6D;
  assign str_print[1184] = 8'h5F;
  assign str_print[1185] = 8'h77;
  assign str_print[1186] = 8'h65;
  assign str_print[1187] = 8'h6E;
  assign str_print[1188] = 8'h3A;
  assign str_print[1189] = 8'h20;
  assign str_print[1191] = 8'h09;
  assign str_print[1192] = 8'h6D;
  assign str_print[1193] = 8'h65;
  assign str_print[1194] = 8'h6D;
  assign str_print[1195] = 8'h5F;
  assign str_print[1196] = 8'h72;
  assign str_print[1197] = 8'h65;
  assign str_print[1198] = 8'h6E;
  assign str_print[1199] = 8'h3A;
  assign str_print[1200] = 8'h20;
  assign str_print[1202] = 8'h09;
  assign str_print[1203] = 8'h69;
  assign str_print[1204] = 8'h73;
  assign str_print[1205] = 8'h5F;
  assign str_print[1206] = 8'h6A;
  assign str_print[1207] = 8'h61;
  assign str_print[1208] = 8'h6C;
  assign str_print[1209] = 8'h3A;
  assign str_print[1210] = 8'h20;
  assign str_print[1212] = 8'h09;
  assign str_print[1213] = 8'h69;
  assign str_print[1214] = 8'h73;
  assign str_print[1215] = 8'h5F;
  assign str_print[1216] = 8'h6A;
  assign str_print[1217] = 8'h61;
  assign str_print[1218] = 8'h6C;
  assign str_print[1219] = 8'h72;
  assign str_print[1220] = 8'h3A;
  assign str_print[1221] = 8'h20;
  assign str_print[1223] = 8'h0A;
  assign str_print[1224] = 8'h0D;
  assign str_print[1225] = 8'h3D;
  assign str_print[1226] = 8'h3D;
  assign str_print[1227] = 8'h3D;
  assign str_print[1228] = 8'h3D;
  assign str_print[1229] = 8'h3D;
  assign str_print[1230] = 8'h3D;
  assign str_print[1231] = 8'h3D;
  assign str_print[1232] = 8'h3D;
  assign str_print[1233] = 8'h3D;
  assign str_print[1234] = 8'h3D;
  assign str_print[1235] = 8'h3D;
  assign str_print[1236] = 8'h3D;
  assign str_print[1237] = 8'h3D;
  assign str_print[1238] = 8'h3D;
  assign str_print[1239] = 8'h3D;
  assign str_print[1240] = 8'h3D;
  assign str_print[1241] = 8'h3D;
  assign str_print[1242] = 8'h3D;
  assign str_print[1243] = 8'h3D;
  assign str_print[1244] = 8'h3D;
  assign str_print[1245] = 8'h3D;
  assign str_print[1246] = 8'h3D;
  assign str_print[1247] = 8'h3D;
  assign str_print[1248] = 8'h3D;
  assign str_print[1249] = 8'h3D;
  assign str_print[1250] = 8'h3D;
  assign str_print[1251] = 8'h3D;
  assign str_print[1252] = 8'h3D;
  assign str_print[1253] = 8'h3D;
  assign str_print[1254] = 8'h3D;
  assign str_print[1255] = 8'h3D;
  assign str_print[1256] = 8'h3D;
  assign str_print[1257] = 8'h3D;
  assign str_print[1258] = 8'h3D;
  assign str_print[1259] = 8'h3D;
  assign str_print[1260] = 8'h3D;
  assign str_print[1261] = 8'h3D;
  assign str_print[1262] = 8'h3D;
  assign str_print[1263] = 8'h20;
  assign str_print[1264] = 8'h57;
  assign str_print[1265] = 8'h62;
  assign str_print[1266] = 8'h20;
  assign str_print[1267] = 8'h3D;
  assign str_print[1268] = 8'h3D;
  assign str_print[1269] = 8'h3D;
  assign str_print[1270] = 8'h3D;
  assign str_print[1271] = 8'h3D;
  assign str_print[1272] = 8'h3D;
  assign str_print[1273] = 8'h3D;
  assign str_print[1274] = 8'h3D;
  assign str_print[1275] = 8'h3D;
  assign str_print[1276] = 8'h3D;
  assign str_print[1277] = 8'h3D;
  assign str_print[1278] = 8'h3D;
  assign str_print[1279] = 8'h3D;
  assign str_print[1280] = 8'h3D;
  assign str_print[1281] = 8'h3D;
  assign str_print[1282] = 8'h3D;
  assign str_print[1283] = 8'h3D;
  assign str_print[1284] = 8'h3D;
  assign str_print[1285] = 8'h3D;
  assign str_print[1286] = 8'h3D;
  assign str_print[1287] = 8'h3D;
  assign str_print[1288] = 8'h3D;
  assign str_print[1289] = 8'h3D;
  assign str_print[1290] = 8'h3D;
  assign str_print[1291] = 8'h3D;
  assign str_print[1292] = 8'h3D;
  assign str_print[1293] = 8'h3D;
  assign str_print[1294] = 8'h3D;
  assign str_print[1295] = 8'h3D;
  assign str_print[1296] = 8'h3D;
  assign str_print[1297] = 8'h3D;
  assign str_print[1298] = 8'h3D;
  assign str_print[1299] = 8'h3D;
  assign str_print[1300] = 8'h3D;
  assign str_print[1301] = 8'h3D;
  assign str_print[1302] = 8'h3D;
  assign str_print[1303] = 8'h3D;
  assign str_print[1304] = 8'h3D;
  assign str_print[1305] = 8'h3D;
  assign str_print[1306] = 8'h0A;
  assign str_print[1307] = 8'h0D;
  assign str_print[1308] = 8'h70;
  assign str_print[1309] = 8'h63;
  assign str_print[1310] = 8'h3A;
  assign str_print[1311] = 8'h20;
  assign str_print[1320] = 8'h09;
  assign str_print[1321] = 8'h69;
  assign str_print[1322] = 8'h6E;
  assign str_print[1323] = 8'h73;
  assign str_print[1324] = 8'h74;
  assign str_print[1325] = 8'h3A;
  assign str_print[1326] = 8'h20;
  assign str_print[1335] = 8'h09;
  assign str_print[1336] = 8'h76;
  assign str_print[1337] = 8'h61;
  assign str_print[1338] = 8'h6C;
  assign str_print[1339] = 8'h69;
  assign str_print[1340] = 8'h64;
  assign str_print[1341] = 8'h3A;
  assign str_print[1342] = 8'h20;
  assign str_print[1344] = 8'h0A;
  assign str_print[1345] = 8'h0D;
  assign str_print[1346] = 8'h72;
  assign str_print[1347] = 8'h64;
  assign str_print[1348] = 8'h3A;
  assign str_print[1349] = 8'h20;
  assign str_print[1350] = 8'h20;
  assign str_print[1353] = 8'h09;
  assign str_print[1354] = 8'h72;
  assign str_print[1355] = 8'h65;
  assign str_print[1356] = 8'h67;
  assign str_print[1357] = 8'h5F;
  assign str_print[1358] = 8'h77;
  assign str_print[1359] = 8'h65;
  assign str_print[1360] = 8'h6E;
  assign str_print[1361] = 8'h3A;
  assign str_print[1362] = 8'h20;
  assign str_print[1364] = 8'h09;
  assign str_print[1365] = 8'h72;
  assign str_print[1366] = 8'h65;
  assign str_print[1367] = 8'h67;
  assign str_print[1368] = 8'h5F;
  assign str_print[1369] = 8'h77;
  assign str_print[1370] = 8'h5F;
  assign str_print[1371] = 8'h64;
  assign str_print[1372] = 8'h61;
  assign str_print[1373] = 8'h74;
  assign str_print[1374] = 8'h61;
  assign str_print[1375] = 8'h3A;
  assign str_print[1376] = 8'h20;
  assign str_print[1385] = 8'h0D;
  assign str_print[1386] = 8'h08;
  assign str_print[1387] = 8'h0D;
  assign str_print[1388] = 8'h08;
  assign str_print[1389] = 8'h0D;
  assign str_print[1390] = 8'h08;
  assign str_print[1391] = 8'h0D;
  assign str_print[1392] = 8'h08;
  assign str_print[1393] = 8'h0D;
  assign str_print[1394] = 8'h08;
  assign str_print[1395] = 8'h0D;
  assign str_print[1396] = 8'h08;
  assign str_print[1397] = 8'h0D;
  assign str_print[1398] = 8'h08;
  assign str_print[1399] = 8'h0D;
  assign str_print[1400] = 8'h08;
  assign str_print[1401] = 8'h0D;
  assign str_print[1402] = 8'h08;
  assign str_print[1403] = 8'h0D;
  assign str_print[1404] = 8'h08;
  assign str_print[1405] = 8'h0D;
  assign str_print[1406] = 8'h08;
  assign str_print[1407] = 8'h0D;
  assign str_print[1408] = 8'h08;
  assign str_print[1409] = 8'h0D;
  assign str_print[1410] = 8'h08;
  assign str_print[1411] = 8'h0D;
  assign str_print[1412] = 8'h08;
  assign str_print[1413] = 8'h0D;
  assign str_print[1414] = 8'h08;
  assign str_print[1415] = 8'h0D;
  assign str_print[1416] = 8'h08;
  assign str_print[1417] = 8'h0D;
  assign str_print[1418] = 8'h08;
  assign str_print[1419] = 8'h0D;
  assign str_print[1420] = 8'h08;
  assign str_print[1421] = 8'h0D;
  assign str_print[1422] = 8'h08;
  assign str_print[1423] = 8'h0D;
  assign str_print[1424] = 8'h08;
  assign str_print[1425] = 8'h0D;
  assign str_print[1426] = 8'h08;
  assign str_print[1427] = 8'h0D;
  assign str_print[1428] = 8'h08;
  assign str_print[1429] = 8'h0D;
  assign str_print[1430] = 8'h08;
  assign str_print[1431] = 8'h0D;
  assign str_print[1432] = 8'h08;
  assign str_print[1433] = 8'h0D;
  assign str_print[1434] = 8'h08;
  assign str_print[1435] = 8'h0D;


  // Instance for hex2ascii
  hex_to_ascii inst_pc_if_7 (.hex(pc_if[31:28]), .ascii(str_print[110]));
  hex_to_ascii inst_pc_if_6 (.hex(pc_if[27:24]), .ascii(str_print[111]));
  hex_to_ascii inst_pc_if_5 (.hex(pc_if[23:20]), .ascii(str_print[112]));
  hex_to_ascii inst_pc_if_4 (.hex(pc_if[19:16]), .ascii(str_print[113]));
  hex_to_ascii inst_pc_if_3 (.hex(pc_if[15:12]), .ascii(str_print[114]));
  hex_to_ascii inst_pc_if_2 (.hex(pc_if[11:8]), .ascii(str_print[115]));
  hex_to_ascii inst_pc_if_1 (.hex(pc_if[7:4]), .ascii(str_print[116]));
  hex_to_ascii inst_pc_if_0 (.hex(pc_if[3:0]), .ascii(str_print[117]));
  hex_to_ascii inst_inst_if_7 (.hex(inst_if[31:28]), .ascii(str_print[125]));
  hex_to_ascii inst_inst_if_6 (.hex(inst_if[27:24]), .ascii(str_print[126]));
  hex_to_ascii inst_inst_if_5 (.hex(inst_if[23:20]), .ascii(str_print[127]));
  hex_to_ascii inst_inst_if_4 (.hex(inst_if[19:16]), .ascii(str_print[128]));
  hex_to_ascii inst_inst_if_3 (.hex(inst_if[15:12]), .ascii(str_print[129]));
  hex_to_ascii inst_inst_if_2 (.hex(inst_if[11:8]), .ascii(str_print[130]));
  hex_to_ascii inst_inst_if_1 (.hex(inst_if[7:4]), .ascii(str_print[131]));
  hex_to_ascii inst_inst_if_0 (.hex(inst_if[3:0]), .ascii(str_print[132]));
  hex_to_ascii inst_pc_id_7 (.hex(pc_id[31:28]), .ascii(str_print[222]));
  hex_to_ascii inst_pc_id_6 (.hex(pc_id[27:24]), .ascii(str_print[223]));
  hex_to_ascii inst_pc_id_5 (.hex(pc_id[23:20]), .ascii(str_print[224]));
  hex_to_ascii inst_pc_id_4 (.hex(pc_id[19:16]), .ascii(str_print[225]));
  hex_to_ascii inst_pc_id_3 (.hex(pc_id[15:12]), .ascii(str_print[226]));
  hex_to_ascii inst_pc_id_2 (.hex(pc_id[11:8]), .ascii(str_print[227]));
  hex_to_ascii inst_pc_id_1 (.hex(pc_id[7:4]), .ascii(str_print[228]));
  hex_to_ascii inst_pc_id_0 (.hex(pc_id[3:0]), .ascii(str_print[229]));
  hex_to_ascii inst_inst_id_7 (.hex(inst_id[31:28]), .ascii(str_print[237]));
  hex_to_ascii inst_inst_id_6 (.hex(inst_id[27:24]), .ascii(str_print[238]));
  hex_to_ascii inst_inst_id_5 (.hex(inst_id[23:20]), .ascii(str_print[239]));
  hex_to_ascii inst_inst_id_4 (.hex(inst_id[19:16]), .ascii(str_print[240]));
  hex_to_ascii inst_inst_id_3 (.hex(inst_id[15:12]), .ascii(str_print[241]));
  hex_to_ascii inst_inst_id_2 (.hex(inst_id[11:8]), .ascii(str_print[242]));
  hex_to_ascii inst_inst_id_1 (.hex(inst_id[7:4]), .ascii(str_print[243]));
  hex_to_ascii inst_inst_id_0 (.hex(inst_id[3:0]), .ascii(str_print[244]));
  hex_to_ascii inst_valid_id_0 (.hex({3'b0,valid_id}), .ascii(str_print[253]));
  hex_to_ascii inst_x0_7 (.hex(x0[31:28]), .ascii(str_print[260]));
  hex_to_ascii inst_x0_6 (.hex(x0[27:24]), .ascii(str_print[261]));
  hex_to_ascii inst_x0_5 (.hex(x0[23:20]), .ascii(str_print[262]));
  hex_to_ascii inst_x0_4 (.hex(x0[19:16]), .ascii(str_print[263]));
  hex_to_ascii inst_x0_3 (.hex(x0[15:12]), .ascii(str_print[264]));
  hex_to_ascii inst_x0_2 (.hex(x0[11:8]), .ascii(str_print[265]));
  hex_to_ascii inst_x0_1 (.hex(x0[7:4]), .ascii(str_print[266]));
  hex_to_ascii inst_x0_0 (.hex(x0[3:0]), .ascii(str_print[267]));
  hex_to_ascii inst_ra_7 (.hex(ra[31:28]), .ascii(str_print[273]));
  hex_to_ascii inst_ra_6 (.hex(ra[27:24]), .ascii(str_print[274]));
  hex_to_ascii inst_ra_5 (.hex(ra[23:20]), .ascii(str_print[275]));
  hex_to_ascii inst_ra_4 (.hex(ra[19:16]), .ascii(str_print[276]));
  hex_to_ascii inst_ra_3 (.hex(ra[15:12]), .ascii(str_print[277]));
  hex_to_ascii inst_ra_2 (.hex(ra[11:8]), .ascii(str_print[278]));
  hex_to_ascii inst_ra_1 (.hex(ra[7:4]), .ascii(str_print[279]));
  hex_to_ascii inst_ra_0 (.hex(ra[3:0]), .ascii(str_print[280]));
  hex_to_ascii inst_sp_7 (.hex(sp[31:28]), .ascii(str_print[286]));
  hex_to_ascii inst_sp_6 (.hex(sp[27:24]), .ascii(str_print[287]));
  hex_to_ascii inst_sp_5 (.hex(sp[23:20]), .ascii(str_print[288]));
  hex_to_ascii inst_sp_4 (.hex(sp[19:16]), .ascii(str_print[289]));
  hex_to_ascii inst_sp_3 (.hex(sp[15:12]), .ascii(str_print[290]));
  hex_to_ascii inst_sp_2 (.hex(sp[11:8]), .ascii(str_print[291]));
  hex_to_ascii inst_sp_1 (.hex(sp[7:4]), .ascii(str_print[292]));
  hex_to_ascii inst_sp_0 (.hex(sp[3:0]), .ascii(str_print[293]));
  hex_to_ascii inst_gp_7 (.hex(gp[31:28]), .ascii(str_print[299]));
  hex_to_ascii inst_gp_6 (.hex(gp[27:24]), .ascii(str_print[300]));
  hex_to_ascii inst_gp_5 (.hex(gp[23:20]), .ascii(str_print[301]));
  hex_to_ascii inst_gp_4 (.hex(gp[19:16]), .ascii(str_print[302]));
  hex_to_ascii inst_gp_3 (.hex(gp[15:12]), .ascii(str_print[303]));
  hex_to_ascii inst_gp_2 (.hex(gp[11:8]), .ascii(str_print[304]));
  hex_to_ascii inst_gp_1 (.hex(gp[7:4]), .ascii(str_print[305]));
  hex_to_ascii inst_gp_0 (.hex(gp[3:0]), .ascii(str_print[306]));
  hex_to_ascii inst_tp_7 (.hex(tp[31:28]), .ascii(str_print[312]));
  hex_to_ascii inst_tp_6 (.hex(tp[27:24]), .ascii(str_print[313]));
  hex_to_ascii inst_tp_5 (.hex(tp[23:20]), .ascii(str_print[314]));
  hex_to_ascii inst_tp_4 (.hex(tp[19:16]), .ascii(str_print[315]));
  hex_to_ascii inst_tp_3 (.hex(tp[15:12]), .ascii(str_print[316]));
  hex_to_ascii inst_tp_2 (.hex(tp[11:8]), .ascii(str_print[317]));
  hex_to_ascii inst_tp_1 (.hex(tp[7:4]), .ascii(str_print[318]));
  hex_to_ascii inst_tp_0 (.hex(tp[3:0]), .ascii(str_print[319]));
  hex_to_ascii inst_t0_7 (.hex(t0[31:28]), .ascii(str_print[326]));
  hex_to_ascii inst_t0_6 (.hex(t0[27:24]), .ascii(str_print[327]));
  hex_to_ascii inst_t0_5 (.hex(t0[23:20]), .ascii(str_print[328]));
  hex_to_ascii inst_t0_4 (.hex(t0[19:16]), .ascii(str_print[329]));
  hex_to_ascii inst_t0_3 (.hex(t0[15:12]), .ascii(str_print[330]));
  hex_to_ascii inst_t0_2 (.hex(t0[11:8]), .ascii(str_print[331]));
  hex_to_ascii inst_t0_1 (.hex(t0[7:4]), .ascii(str_print[332]));
  hex_to_ascii inst_t0_0 (.hex(t0[3:0]), .ascii(str_print[333]));
  hex_to_ascii inst_t1_7 (.hex(t1[31:28]), .ascii(str_print[339]));
  hex_to_ascii inst_t1_6 (.hex(t1[27:24]), .ascii(str_print[340]));
  hex_to_ascii inst_t1_5 (.hex(t1[23:20]), .ascii(str_print[341]));
  hex_to_ascii inst_t1_4 (.hex(t1[19:16]), .ascii(str_print[342]));
  hex_to_ascii inst_t1_3 (.hex(t1[15:12]), .ascii(str_print[343]));
  hex_to_ascii inst_t1_2 (.hex(t1[11:8]), .ascii(str_print[344]));
  hex_to_ascii inst_t1_1 (.hex(t1[7:4]), .ascii(str_print[345]));
  hex_to_ascii inst_t1_0 (.hex(t1[3:0]), .ascii(str_print[346]));
  hex_to_ascii inst_t2_7 (.hex(t2[31:28]), .ascii(str_print[352]));
  hex_to_ascii inst_t2_6 (.hex(t2[27:24]), .ascii(str_print[353]));
  hex_to_ascii inst_t2_5 (.hex(t2[23:20]), .ascii(str_print[354]));
  hex_to_ascii inst_t2_4 (.hex(t2[19:16]), .ascii(str_print[355]));
  hex_to_ascii inst_t2_3 (.hex(t2[15:12]), .ascii(str_print[356]));
  hex_to_ascii inst_t2_2 (.hex(t2[11:8]), .ascii(str_print[357]));
  hex_to_ascii inst_t2_1 (.hex(t2[7:4]), .ascii(str_print[358]));
  hex_to_ascii inst_t2_0 (.hex(t2[3:0]), .ascii(str_print[359]));
  hex_to_ascii inst_s0_7 (.hex(s0[31:28]), .ascii(str_print[365]));
  hex_to_ascii inst_s0_6 (.hex(s0[27:24]), .ascii(str_print[366]));
  hex_to_ascii inst_s0_5 (.hex(s0[23:20]), .ascii(str_print[367]));
  hex_to_ascii inst_s0_4 (.hex(s0[19:16]), .ascii(str_print[368]));
  hex_to_ascii inst_s0_3 (.hex(s0[15:12]), .ascii(str_print[369]));
  hex_to_ascii inst_s0_2 (.hex(s0[11:8]), .ascii(str_print[370]));
  hex_to_ascii inst_s0_1 (.hex(s0[7:4]), .ascii(str_print[371]));
  hex_to_ascii inst_s0_0 (.hex(s0[3:0]), .ascii(str_print[372]));
  hex_to_ascii inst_s1_7 (.hex(s1[31:28]), .ascii(str_print[378]));
  hex_to_ascii inst_s1_6 (.hex(s1[27:24]), .ascii(str_print[379]));
  hex_to_ascii inst_s1_5 (.hex(s1[23:20]), .ascii(str_print[380]));
  hex_to_ascii inst_s1_4 (.hex(s1[19:16]), .ascii(str_print[381]));
  hex_to_ascii inst_s1_3 (.hex(s1[15:12]), .ascii(str_print[382]));
  hex_to_ascii inst_s1_2 (.hex(s1[11:8]), .ascii(str_print[383]));
  hex_to_ascii inst_s1_1 (.hex(s1[7:4]), .ascii(str_print[384]));
  hex_to_ascii inst_s1_0 (.hex(s1[3:0]), .ascii(str_print[385]));
  hex_to_ascii inst_a0_7 (.hex(a0[31:28]), .ascii(str_print[392]));
  hex_to_ascii inst_a0_6 (.hex(a0[27:24]), .ascii(str_print[393]));
  hex_to_ascii inst_a0_5 (.hex(a0[23:20]), .ascii(str_print[394]));
  hex_to_ascii inst_a0_4 (.hex(a0[19:16]), .ascii(str_print[395]));
  hex_to_ascii inst_a0_3 (.hex(a0[15:12]), .ascii(str_print[396]));
  hex_to_ascii inst_a0_2 (.hex(a0[11:8]), .ascii(str_print[397]));
  hex_to_ascii inst_a0_1 (.hex(a0[7:4]), .ascii(str_print[398]));
  hex_to_ascii inst_a0_0 (.hex(a0[3:0]), .ascii(str_print[399]));
  hex_to_ascii inst_a1_7 (.hex(a1[31:28]), .ascii(str_print[405]));
  hex_to_ascii inst_a1_6 (.hex(a1[27:24]), .ascii(str_print[406]));
  hex_to_ascii inst_a1_5 (.hex(a1[23:20]), .ascii(str_print[407]));
  hex_to_ascii inst_a1_4 (.hex(a1[19:16]), .ascii(str_print[408]));
  hex_to_ascii inst_a1_3 (.hex(a1[15:12]), .ascii(str_print[409]));
  hex_to_ascii inst_a1_2 (.hex(a1[11:8]), .ascii(str_print[410]));
  hex_to_ascii inst_a1_1 (.hex(a1[7:4]), .ascii(str_print[411]));
  hex_to_ascii inst_a1_0 (.hex(a1[3:0]), .ascii(str_print[412]));
  hex_to_ascii inst_a2_7 (.hex(a2[31:28]), .ascii(str_print[418]));
  hex_to_ascii inst_a2_6 (.hex(a2[27:24]), .ascii(str_print[419]));
  hex_to_ascii inst_a2_5 (.hex(a2[23:20]), .ascii(str_print[420]));
  hex_to_ascii inst_a2_4 (.hex(a2[19:16]), .ascii(str_print[421]));
  hex_to_ascii inst_a2_3 (.hex(a2[15:12]), .ascii(str_print[422]));
  hex_to_ascii inst_a2_2 (.hex(a2[11:8]), .ascii(str_print[423]));
  hex_to_ascii inst_a2_1 (.hex(a2[7:4]), .ascii(str_print[424]));
  hex_to_ascii inst_a2_0 (.hex(a2[3:0]), .ascii(str_print[425]));
  hex_to_ascii inst_a3_7 (.hex(a3[31:28]), .ascii(str_print[431]));
  hex_to_ascii inst_a3_6 (.hex(a3[27:24]), .ascii(str_print[432]));
  hex_to_ascii inst_a3_5 (.hex(a3[23:20]), .ascii(str_print[433]));
  hex_to_ascii inst_a3_4 (.hex(a3[19:16]), .ascii(str_print[434]));
  hex_to_ascii inst_a3_3 (.hex(a3[15:12]), .ascii(str_print[435]));
  hex_to_ascii inst_a3_2 (.hex(a3[11:8]), .ascii(str_print[436]));
  hex_to_ascii inst_a3_1 (.hex(a3[7:4]), .ascii(str_print[437]));
  hex_to_ascii inst_a3_0 (.hex(a3[3:0]), .ascii(str_print[438]));
  hex_to_ascii inst_a4_7 (.hex(a4[31:28]), .ascii(str_print[444]));
  hex_to_ascii inst_a4_6 (.hex(a4[27:24]), .ascii(str_print[445]));
  hex_to_ascii inst_a4_5 (.hex(a4[23:20]), .ascii(str_print[446]));
  hex_to_ascii inst_a4_4 (.hex(a4[19:16]), .ascii(str_print[447]));
  hex_to_ascii inst_a4_3 (.hex(a4[15:12]), .ascii(str_print[448]));
  hex_to_ascii inst_a4_2 (.hex(a4[11:8]), .ascii(str_print[449]));
  hex_to_ascii inst_a4_1 (.hex(a4[7:4]), .ascii(str_print[450]));
  hex_to_ascii inst_a4_0 (.hex(a4[3:0]), .ascii(str_print[451]));
  hex_to_ascii inst_a5_7 (.hex(a5[31:28]), .ascii(str_print[458]));
  hex_to_ascii inst_a5_6 (.hex(a5[27:24]), .ascii(str_print[459]));
  hex_to_ascii inst_a5_5 (.hex(a5[23:20]), .ascii(str_print[460]));
  hex_to_ascii inst_a5_4 (.hex(a5[19:16]), .ascii(str_print[461]));
  hex_to_ascii inst_a5_3 (.hex(a5[15:12]), .ascii(str_print[462]));
  hex_to_ascii inst_a5_2 (.hex(a5[11:8]), .ascii(str_print[463]));
  hex_to_ascii inst_a5_1 (.hex(a5[7:4]), .ascii(str_print[464]));
  hex_to_ascii inst_a5_0 (.hex(a5[3:0]), .ascii(str_print[465]));
  hex_to_ascii inst_a6_7 (.hex(a6[31:28]), .ascii(str_print[471]));
  hex_to_ascii inst_a6_6 (.hex(a6[27:24]), .ascii(str_print[472]));
  hex_to_ascii inst_a6_5 (.hex(a6[23:20]), .ascii(str_print[473]));
  hex_to_ascii inst_a6_4 (.hex(a6[19:16]), .ascii(str_print[474]));
  hex_to_ascii inst_a6_3 (.hex(a6[15:12]), .ascii(str_print[475]));
  hex_to_ascii inst_a6_2 (.hex(a6[11:8]), .ascii(str_print[476]));
  hex_to_ascii inst_a6_1 (.hex(a6[7:4]), .ascii(str_print[477]));
  hex_to_ascii inst_a6_0 (.hex(a6[3:0]), .ascii(str_print[478]));
  hex_to_ascii inst_a7_7 (.hex(a7[31:28]), .ascii(str_print[484]));
  hex_to_ascii inst_a7_6 (.hex(a7[27:24]), .ascii(str_print[485]));
  hex_to_ascii inst_a7_5 (.hex(a7[23:20]), .ascii(str_print[486]));
  hex_to_ascii inst_a7_4 (.hex(a7[19:16]), .ascii(str_print[487]));
  hex_to_ascii inst_a7_3 (.hex(a7[15:12]), .ascii(str_print[488]));
  hex_to_ascii inst_a7_2 (.hex(a7[11:8]), .ascii(str_print[489]));
  hex_to_ascii inst_a7_1 (.hex(a7[7:4]), .ascii(str_print[490]));
  hex_to_ascii inst_a7_0 (.hex(a7[3:0]), .ascii(str_print[491]));
  hex_to_ascii inst_s2_7 (.hex(s2[31:28]), .ascii(str_print[497]));
  hex_to_ascii inst_s2_6 (.hex(s2[27:24]), .ascii(str_print[498]));
  hex_to_ascii inst_s2_5 (.hex(s2[23:20]), .ascii(str_print[499]));
  hex_to_ascii inst_s2_4 (.hex(s2[19:16]), .ascii(str_print[500]));
  hex_to_ascii inst_s2_3 (.hex(s2[15:12]), .ascii(str_print[501]));
  hex_to_ascii inst_s2_2 (.hex(s2[11:8]), .ascii(str_print[502]));
  hex_to_ascii inst_s2_1 (.hex(s2[7:4]), .ascii(str_print[503]));
  hex_to_ascii inst_s2_0 (.hex(s2[3:0]), .ascii(str_print[504]));
  hex_to_ascii inst_s3_7 (.hex(s3[31:28]), .ascii(str_print[510]));
  hex_to_ascii inst_s3_6 (.hex(s3[27:24]), .ascii(str_print[511]));
  hex_to_ascii inst_s3_5 (.hex(s3[23:20]), .ascii(str_print[512]));
  hex_to_ascii inst_s3_4 (.hex(s3[19:16]), .ascii(str_print[513]));
  hex_to_ascii inst_s3_3 (.hex(s3[15:12]), .ascii(str_print[514]));
  hex_to_ascii inst_s3_2 (.hex(s3[11:8]), .ascii(str_print[515]));
  hex_to_ascii inst_s3_1 (.hex(s3[7:4]), .ascii(str_print[516]));
  hex_to_ascii inst_s3_0 (.hex(s3[3:0]), .ascii(str_print[517]));
  hex_to_ascii inst_s4_7 (.hex(s4[31:28]), .ascii(str_print[524]));
  hex_to_ascii inst_s4_6 (.hex(s4[27:24]), .ascii(str_print[525]));
  hex_to_ascii inst_s4_5 (.hex(s4[23:20]), .ascii(str_print[526]));
  hex_to_ascii inst_s4_4 (.hex(s4[19:16]), .ascii(str_print[527]));
  hex_to_ascii inst_s4_3 (.hex(s4[15:12]), .ascii(str_print[528]));
  hex_to_ascii inst_s4_2 (.hex(s4[11:8]), .ascii(str_print[529]));
  hex_to_ascii inst_s4_1 (.hex(s4[7:4]), .ascii(str_print[530]));
  hex_to_ascii inst_s4_0 (.hex(s4[3:0]), .ascii(str_print[531]));
  hex_to_ascii inst_s5_7 (.hex(s5[31:28]), .ascii(str_print[537]));
  hex_to_ascii inst_s5_6 (.hex(s5[27:24]), .ascii(str_print[538]));
  hex_to_ascii inst_s5_5 (.hex(s5[23:20]), .ascii(str_print[539]));
  hex_to_ascii inst_s5_4 (.hex(s5[19:16]), .ascii(str_print[540]));
  hex_to_ascii inst_s5_3 (.hex(s5[15:12]), .ascii(str_print[541]));
  hex_to_ascii inst_s5_2 (.hex(s5[11:8]), .ascii(str_print[542]));
  hex_to_ascii inst_s5_1 (.hex(s5[7:4]), .ascii(str_print[543]));
  hex_to_ascii inst_s5_0 (.hex(s5[3:0]), .ascii(str_print[544]));
  hex_to_ascii inst_s6_7 (.hex(s6[31:28]), .ascii(str_print[550]));
  hex_to_ascii inst_s6_6 (.hex(s6[27:24]), .ascii(str_print[551]));
  hex_to_ascii inst_s6_5 (.hex(s6[23:20]), .ascii(str_print[552]));
  hex_to_ascii inst_s6_4 (.hex(s6[19:16]), .ascii(str_print[553]));
  hex_to_ascii inst_s6_3 (.hex(s6[15:12]), .ascii(str_print[554]));
  hex_to_ascii inst_s6_2 (.hex(s6[11:8]), .ascii(str_print[555]));
  hex_to_ascii inst_s6_1 (.hex(s6[7:4]), .ascii(str_print[556]));
  hex_to_ascii inst_s6_0 (.hex(s6[3:0]), .ascii(str_print[557]));
  hex_to_ascii inst_s7_7 (.hex(s7[31:28]), .ascii(str_print[563]));
  hex_to_ascii inst_s7_6 (.hex(s7[27:24]), .ascii(str_print[564]));
  hex_to_ascii inst_s7_5 (.hex(s7[23:20]), .ascii(str_print[565]));
  hex_to_ascii inst_s7_4 (.hex(s7[19:16]), .ascii(str_print[566]));
  hex_to_ascii inst_s7_3 (.hex(s7[15:12]), .ascii(str_print[567]));
  hex_to_ascii inst_s7_2 (.hex(s7[11:8]), .ascii(str_print[568]));
  hex_to_ascii inst_s7_1 (.hex(s7[7:4]), .ascii(str_print[569]));
  hex_to_ascii inst_s7_0 (.hex(s7[3:0]), .ascii(str_print[570]));
  hex_to_ascii inst_s8_7 (.hex(s8[31:28]), .ascii(str_print[576]));
  hex_to_ascii inst_s8_6 (.hex(s8[27:24]), .ascii(str_print[577]));
  hex_to_ascii inst_s8_5 (.hex(s8[23:20]), .ascii(str_print[578]));
  hex_to_ascii inst_s8_4 (.hex(s8[19:16]), .ascii(str_print[579]));
  hex_to_ascii inst_s8_3 (.hex(s8[15:12]), .ascii(str_print[580]));
  hex_to_ascii inst_s8_2 (.hex(s8[11:8]), .ascii(str_print[581]));
  hex_to_ascii inst_s8_1 (.hex(s8[7:4]), .ascii(str_print[582]));
  hex_to_ascii inst_s8_0 (.hex(s8[3:0]), .ascii(str_print[583]));
  hex_to_ascii inst_s9_7 (.hex(s9[31:28]), .ascii(str_print[590]));
  hex_to_ascii inst_s9_6 (.hex(s9[27:24]), .ascii(str_print[591]));
  hex_to_ascii inst_s9_5 (.hex(s9[23:20]), .ascii(str_print[592]));
  hex_to_ascii inst_s9_4 (.hex(s9[19:16]), .ascii(str_print[593]));
  hex_to_ascii inst_s9_3 (.hex(s9[15:12]), .ascii(str_print[594]));
  hex_to_ascii inst_s9_2 (.hex(s9[11:8]), .ascii(str_print[595]));
  hex_to_ascii inst_s9_1 (.hex(s9[7:4]), .ascii(str_print[596]));
  hex_to_ascii inst_s9_0 (.hex(s9[3:0]), .ascii(str_print[597]));
  hex_to_ascii inst_s10_7 (.hex(s10[31:28]), .ascii(str_print[603]));
  hex_to_ascii inst_s10_6 (.hex(s10[27:24]), .ascii(str_print[604]));
  hex_to_ascii inst_s10_5 (.hex(s10[23:20]), .ascii(str_print[605]));
  hex_to_ascii inst_s10_4 (.hex(s10[19:16]), .ascii(str_print[606]));
  hex_to_ascii inst_s10_3 (.hex(s10[15:12]), .ascii(str_print[607]));
  hex_to_ascii inst_s10_2 (.hex(s10[11:8]), .ascii(str_print[608]));
  hex_to_ascii inst_s10_1 (.hex(s10[7:4]), .ascii(str_print[609]));
  hex_to_ascii inst_s10_0 (.hex(s10[3:0]), .ascii(str_print[610]));
  hex_to_ascii inst_s11_7 (.hex(s11[31:28]), .ascii(str_print[616]));
  hex_to_ascii inst_s11_6 (.hex(s11[27:24]), .ascii(str_print[617]));
  hex_to_ascii inst_s11_5 (.hex(s11[23:20]), .ascii(str_print[618]));
  hex_to_ascii inst_s11_4 (.hex(s11[19:16]), .ascii(str_print[619]));
  hex_to_ascii inst_s11_3 (.hex(s11[15:12]), .ascii(str_print[620]));
  hex_to_ascii inst_s11_2 (.hex(s11[11:8]), .ascii(str_print[621]));
  hex_to_ascii inst_s11_1 (.hex(s11[7:4]), .ascii(str_print[622]));
  hex_to_ascii inst_s11_0 (.hex(s11[3:0]), .ascii(str_print[623]));
  hex_to_ascii inst_t3_7 (.hex(t3[31:28]), .ascii(str_print[629]));
  hex_to_ascii inst_t3_6 (.hex(t3[27:24]), .ascii(str_print[630]));
  hex_to_ascii inst_t3_5 (.hex(t3[23:20]), .ascii(str_print[631]));
  hex_to_ascii inst_t3_4 (.hex(t3[19:16]), .ascii(str_print[632]));
  hex_to_ascii inst_t3_3 (.hex(t3[15:12]), .ascii(str_print[633]));
  hex_to_ascii inst_t3_2 (.hex(t3[11:8]), .ascii(str_print[634]));
  hex_to_ascii inst_t3_1 (.hex(t3[7:4]), .ascii(str_print[635]));
  hex_to_ascii inst_t3_0 (.hex(t3[3:0]), .ascii(str_print[636]));
  hex_to_ascii inst_t4_7 (.hex(t4[31:28]), .ascii(str_print[642]));
  hex_to_ascii inst_t4_6 (.hex(t4[27:24]), .ascii(str_print[643]));
  hex_to_ascii inst_t4_5 (.hex(t4[23:20]), .ascii(str_print[644]));
  hex_to_ascii inst_t4_4 (.hex(t4[19:16]), .ascii(str_print[645]));
  hex_to_ascii inst_t4_3 (.hex(t4[15:12]), .ascii(str_print[646]));
  hex_to_ascii inst_t4_2 (.hex(t4[11:8]), .ascii(str_print[647]));
  hex_to_ascii inst_t4_1 (.hex(t4[7:4]), .ascii(str_print[648]));
  hex_to_ascii inst_t4_0 (.hex(t4[3:0]), .ascii(str_print[649]));
  hex_to_ascii inst_t5_7 (.hex(t5[31:28]), .ascii(str_print[656]));
  hex_to_ascii inst_t5_6 (.hex(t5[27:24]), .ascii(str_print[657]));
  hex_to_ascii inst_t5_5 (.hex(t5[23:20]), .ascii(str_print[658]));
  hex_to_ascii inst_t5_4 (.hex(t5[19:16]), .ascii(str_print[659]));
  hex_to_ascii inst_t5_3 (.hex(t5[15:12]), .ascii(str_print[660]));
  hex_to_ascii inst_t5_2 (.hex(t5[11:8]), .ascii(str_print[661]));
  hex_to_ascii inst_t5_1 (.hex(t5[7:4]), .ascii(str_print[662]));
  hex_to_ascii inst_t5_0 (.hex(t5[3:0]), .ascii(str_print[663]));
  hex_to_ascii inst_t6_7 (.hex(t6[31:28]), .ascii(str_print[669]));
  hex_to_ascii inst_t6_6 (.hex(t6[27:24]), .ascii(str_print[670]));
  hex_to_ascii inst_t6_5 (.hex(t6[23:20]), .ascii(str_print[671]));
  hex_to_ascii inst_t6_4 (.hex(t6[19:16]), .ascii(str_print[672]));
  hex_to_ascii inst_t6_3 (.hex(t6[15:12]), .ascii(str_print[673]));
  hex_to_ascii inst_t6_2 (.hex(t6[11:8]), .ascii(str_print[674]));
  hex_to_ascii inst_t6_1 (.hex(t6[7:4]), .ascii(str_print[675]));
  hex_to_ascii inst_t6_0 (.hex(t6[3:0]), .ascii(str_print[676]));
  hex_to_ascii inst_pc_ex_7 (.hex(pc_ex[31:28]), .ascii(str_print[766]));
  hex_to_ascii inst_pc_ex_6 (.hex(pc_ex[27:24]), .ascii(str_print[767]));
  hex_to_ascii inst_pc_ex_5 (.hex(pc_ex[23:20]), .ascii(str_print[768]));
  hex_to_ascii inst_pc_ex_4 (.hex(pc_ex[19:16]), .ascii(str_print[769]));
  hex_to_ascii inst_pc_ex_3 (.hex(pc_ex[15:12]), .ascii(str_print[770]));
  hex_to_ascii inst_pc_ex_2 (.hex(pc_ex[11:8]), .ascii(str_print[771]));
  hex_to_ascii inst_pc_ex_1 (.hex(pc_ex[7:4]), .ascii(str_print[772]));
  hex_to_ascii inst_pc_ex_0 (.hex(pc_ex[3:0]), .ascii(str_print[773]));
  hex_to_ascii inst_inst_ex_7 (.hex(inst_ex[31:28]), .ascii(str_print[781]));
  hex_to_ascii inst_inst_ex_6 (.hex(inst_ex[27:24]), .ascii(str_print[782]));
  hex_to_ascii inst_inst_ex_5 (.hex(inst_ex[23:20]), .ascii(str_print[783]));
  hex_to_ascii inst_inst_ex_4 (.hex(inst_ex[19:16]), .ascii(str_print[784]));
  hex_to_ascii inst_inst_ex_3 (.hex(inst_ex[15:12]), .ascii(str_print[785]));
  hex_to_ascii inst_inst_ex_2 (.hex(inst_ex[11:8]), .ascii(str_print[786]));
  hex_to_ascii inst_inst_ex_1 (.hex(inst_ex[7:4]), .ascii(str_print[787]));
  hex_to_ascii inst_inst_ex_0 (.hex(inst_ex[3:0]), .ascii(str_print[788]));
  hex_to_ascii inst_valid_ex_0 (.hex({3'b0,valid_ex}), .ascii(str_print[797]));
  hex_to_ascii inst_rd_ex_1 (.hex({3'b0,rd_ex[4]}), .ascii(str_print[805]));
  hex_to_ascii inst_rd_ex_0 (.hex(rd_ex[3:0]), .ascii(str_print[806]));
  hex_to_ascii inst_rs1_1 (.hex({3'b0,rs1[4]}), .ascii(str_print[813]));
  hex_to_ascii inst_rs1_0 (.hex(rs1[3:0]), .ascii(str_print[814]));
  hex_to_ascii inst_rs2_1 (.hex({3'b0,rs2[4]}), .ascii(str_print[821]));
  hex_to_ascii inst_rs2_0 (.hex(rs2[3:0]), .ascii(str_print[822]));
  hex_to_ascii inst_rs1_val_7 (.hex(rs1_val[31:28]), .ascii(str_print[833]));
  hex_to_ascii inst_rs1_val_6 (.hex(rs1_val[27:24]), .ascii(str_print[834]));
  hex_to_ascii inst_rs1_val_5 (.hex(rs1_val[23:20]), .ascii(str_print[835]));
  hex_to_ascii inst_rs1_val_4 (.hex(rs1_val[19:16]), .ascii(str_print[836]));
  hex_to_ascii inst_rs1_val_3 (.hex(rs1_val[15:12]), .ascii(str_print[837]));
  hex_to_ascii inst_rs1_val_2 (.hex(rs1_val[11:8]), .ascii(str_print[838]));
  hex_to_ascii inst_rs1_val_1 (.hex(rs1_val[7:4]), .ascii(str_print[839]));
  hex_to_ascii inst_rs1_val_0 (.hex(rs1_val[3:0]), .ascii(str_print[840]));
  hex_to_ascii inst_rs2_val_7 (.hex(rs2_val[31:28]), .ascii(str_print[851]));
  hex_to_ascii inst_rs2_val_6 (.hex(rs2_val[27:24]), .ascii(str_print[852]));
  hex_to_ascii inst_rs2_val_5 (.hex(rs2_val[23:20]), .ascii(str_print[853]));
  hex_to_ascii inst_rs2_val_4 (.hex(rs2_val[19:16]), .ascii(str_print[854]));
  hex_to_ascii inst_rs2_val_3 (.hex(rs2_val[15:12]), .ascii(str_print[855]));
  hex_to_ascii inst_rs2_val_2 (.hex(rs2_val[11:8]), .ascii(str_print[856]));
  hex_to_ascii inst_rs2_val_1 (.hex(rs2_val[7:4]), .ascii(str_print[857]));
  hex_to_ascii inst_rs2_val_0 (.hex(rs2_val[3:0]), .ascii(str_print[858]));
  hex_to_ascii inst_reg_wen_ex_0 (.hex({3'b0,reg_wen_ex}), .ascii(str_print[869]));
  hex_to_ascii inst_is_imm_0 (.hex({3'b0,is_imm}), .ascii(str_print[880]));
  hex_to_ascii inst_imm_7 (.hex(imm[31:28]), .ascii(str_print[887]));
  hex_to_ascii inst_imm_6 (.hex(imm[27:24]), .ascii(str_print[888]));
  hex_to_ascii inst_imm_5 (.hex(imm[23:20]), .ascii(str_print[889]));
  hex_to_ascii inst_imm_4 (.hex(imm[19:16]), .ascii(str_print[890]));
  hex_to_ascii inst_imm_3 (.hex(imm[15:12]), .ascii(str_print[891]));
  hex_to_ascii inst_imm_2 (.hex(imm[11:8]), .ascii(str_print[892]));
  hex_to_ascii inst_imm_1 (.hex(imm[7:4]), .ascii(str_print[893]));
  hex_to_ascii inst_imm_0 (.hex(imm[3:0]), .ascii(str_print[894]));
  hex_to_ascii inst_mem_wen_ex_0 (.hex({3'b0,mem_wen_ex}), .ascii(str_print[906]));
  hex_to_ascii inst_mem_ren_ex_0 (.hex({3'b0,mem_ren_ex}), .ascii(str_print[917]));
  hex_to_ascii inst_is_branch_0 (.hex({3'b0,is_branch}), .ascii(str_print[930]));
  hex_to_ascii inst_is_jal_ex_0 (.hex({3'b0,is_jal_ex}), .ascii(str_print[940]));
  hex_to_ascii inst_is_jalr_ex_0 (.hex({3'b0,is_jalr_ex}), .ascii(str_print[951]));
  hex_to_ascii inst_is_auipc_0 (.hex({3'b0,is_auipc}), .ascii(str_print[964]));
  hex_to_ascii inst_is_lui_0 (.hex({3'b0,is_lui}), .ascii(str_print[974]));
  hex_to_ascii inst_alu_ctrl_0 (.hex(alu_ctrl[3:0]), .ascii(str_print[986]));
  hex_to_ascii inst_cmp_ctrl_0 (.hex({1'b0,cmp_ctrl[2:0]}), .ascii(str_print[998]));
  hex_to_ascii inst_pc_mem_7 (.hex(pc_mem[31:28]), .ascii(str_print[1088]));
  hex_to_ascii inst_pc_mem_6 (.hex(pc_mem[27:24]), .ascii(str_print[1089]));
  hex_to_ascii inst_pc_mem_5 (.hex(pc_mem[23:20]), .ascii(str_print[1090]));
  hex_to_ascii inst_pc_mem_4 (.hex(pc_mem[19:16]), .ascii(str_print[1091]));
  hex_to_ascii inst_pc_mem_3 (.hex(pc_mem[15:12]), .ascii(str_print[1092]));
  hex_to_ascii inst_pc_mem_2 (.hex(pc_mem[11:8]), .ascii(str_print[1093]));
  hex_to_ascii inst_pc_mem_1 (.hex(pc_mem[7:4]), .ascii(str_print[1094]));
  hex_to_ascii inst_pc_mem_0 (.hex(pc_mem[3:0]), .ascii(str_print[1095]));
  hex_to_ascii inst_inst_mem_7 (.hex(inst_mem[31:28]), .ascii(str_print[1103]));
  hex_to_ascii inst_inst_mem_6 (.hex(inst_mem[27:24]), .ascii(str_print[1104]));
  hex_to_ascii inst_inst_mem_5 (.hex(inst_mem[23:20]), .ascii(str_print[1105]));
  hex_to_ascii inst_inst_mem_4 (.hex(inst_mem[19:16]), .ascii(str_print[1106]));
  hex_to_ascii inst_inst_mem_3 (.hex(inst_mem[15:12]), .ascii(str_print[1107]));
  hex_to_ascii inst_inst_mem_2 (.hex(inst_mem[11:8]), .ascii(str_print[1108]));
  hex_to_ascii inst_inst_mem_1 (.hex(inst_mem[7:4]), .ascii(str_print[1109]));
  hex_to_ascii inst_inst_mem_0 (.hex(inst_mem[3:0]), .ascii(str_print[1110]));
  hex_to_ascii inst_valid_mem_0 (.hex({3'b0,valid_mem}), .ascii(str_print[1119]));
  hex_to_ascii inst_rd_mem_1 (.hex({3'b0,rd_mem[4]}), .ascii(str_print[1127]));
  hex_to_ascii inst_rd_mem_0 (.hex(rd_mem[3:0]), .ascii(str_print[1128]));
  hex_to_ascii inst_reg_wen_mem_0 (.hex({3'b0,reg_wen_mem}), .ascii(str_print[1139]));
  hex_to_ascii inst_mem_w_data_7 (.hex(mem_w_data[31:28]), .ascii(str_print[1153]));
  hex_to_ascii inst_mem_w_data_6 (.hex(mem_w_data[27:24]), .ascii(str_print[1154]));
  hex_to_ascii inst_mem_w_data_5 (.hex(mem_w_data[23:20]), .ascii(str_print[1155]));
  hex_to_ascii inst_mem_w_data_4 (.hex(mem_w_data[19:16]), .ascii(str_print[1156]));
  hex_to_ascii inst_mem_w_data_3 (.hex(mem_w_data[15:12]), .ascii(str_print[1157]));
  hex_to_ascii inst_mem_w_data_2 (.hex(mem_w_data[11:8]), .ascii(str_print[1158]));
  hex_to_ascii inst_mem_w_data_1 (.hex(mem_w_data[7:4]), .ascii(str_print[1159]));
  hex_to_ascii inst_mem_w_data_0 (.hex(mem_w_data[3:0]), .ascii(str_print[1160]));
  hex_to_ascii inst_alu_res_7 (.hex(alu_res[31:28]), .ascii(str_print[1171]));
  hex_to_ascii inst_alu_res_6 (.hex(alu_res[27:24]), .ascii(str_print[1172]));
  hex_to_ascii inst_alu_res_5 (.hex(alu_res[23:20]), .ascii(str_print[1173]));
  hex_to_ascii inst_alu_res_4 (.hex(alu_res[19:16]), .ascii(str_print[1174]));
  hex_to_ascii inst_alu_res_3 (.hex(alu_res[15:12]), .ascii(str_print[1175]));
  hex_to_ascii inst_alu_res_2 (.hex(alu_res[11:8]), .ascii(str_print[1176]));
  hex_to_ascii inst_alu_res_1 (.hex(alu_res[7:4]), .ascii(str_print[1177]));
  hex_to_ascii inst_alu_res_0 (.hex(alu_res[3:0]), .ascii(str_print[1178]));
  hex_to_ascii inst_mem_wen_mem_0 (.hex({3'b0,mem_wen_mem}), .ascii(str_print[1190]));
  hex_to_ascii inst_mem_ren_mem_0 (.hex({3'b0,mem_ren_mem}), .ascii(str_print[1201]));
  hex_to_ascii inst_is_jal_mem_0 (.hex({3'b0,is_jal_mem}), .ascii(str_print[1211]));
  hex_to_ascii inst_is_jalr_mem_0 (.hex({3'b0,is_jalr_mem}), .ascii(str_print[1222]));
  hex_to_ascii inst_pc_wb_7 (.hex(pc_wb[31:28]), .ascii(str_print[1312]));
  hex_to_ascii inst_pc_wb_6 (.hex(pc_wb[27:24]), .ascii(str_print[1313]));
  hex_to_ascii inst_pc_wb_5 (.hex(pc_wb[23:20]), .ascii(str_print[1314]));
  hex_to_ascii inst_pc_wb_4 (.hex(pc_wb[19:16]), .ascii(str_print[1315]));
  hex_to_ascii inst_pc_wb_3 (.hex(pc_wb[15:12]), .ascii(str_print[1316]));
  hex_to_ascii inst_pc_wb_2 (.hex(pc_wb[11:8]), .ascii(str_print[1317]));
  hex_to_ascii inst_pc_wb_1 (.hex(pc_wb[7:4]), .ascii(str_print[1318]));
  hex_to_ascii inst_pc_wb_0 (.hex(pc_wb[3:0]), .ascii(str_print[1319]));
  hex_to_ascii inst_inst_wb_7 (.hex(inst_wb[31:28]), .ascii(str_print[1327]));
  hex_to_ascii inst_inst_wb_6 (.hex(inst_wb[27:24]), .ascii(str_print[1328]));
  hex_to_ascii inst_inst_wb_5 (.hex(inst_wb[23:20]), .ascii(str_print[1329]));
  hex_to_ascii inst_inst_wb_4 (.hex(inst_wb[19:16]), .ascii(str_print[1330]));
  hex_to_ascii inst_inst_wb_3 (.hex(inst_wb[15:12]), .ascii(str_print[1331]));
  hex_to_ascii inst_inst_wb_2 (.hex(inst_wb[11:8]), .ascii(str_print[1332]));
  hex_to_ascii inst_inst_wb_1 (.hex(inst_wb[7:4]), .ascii(str_print[1333]));
  hex_to_ascii inst_inst_wb_0 (.hex(inst_wb[3:0]), .ascii(str_print[1334]));
  hex_to_ascii inst_valid_wb_0 (.hex({3'b0,valid_wb}), .ascii(str_print[1343]));
  hex_to_ascii inst_rd_wb_1 (.hex({3'b0,rd_wb[4]}), .ascii(str_print[1351]));
  hex_to_ascii inst_rd_wb_0 (.hex(rd_wb[3:0]), .ascii(str_print[1352]));
  hex_to_ascii inst_reg_wen_wb_0 (.hex({3'b0,reg_wen_wb}), .ascii(str_print[1363]));
  hex_to_ascii inst_reg_w_data_7 (.hex(reg_w_data[31:28]), .ascii(str_print[1377]));
  hex_to_ascii inst_reg_w_data_6 (.hex(reg_w_data[27:24]), .ascii(str_print[1378]));
  hex_to_ascii inst_reg_w_data_5 (.hex(reg_w_data[23:20]), .ascii(str_print[1379]));
  hex_to_ascii inst_reg_w_data_4 (.hex(reg_w_data[19:16]), .ascii(str_print[1380]));
  hex_to_ascii inst_reg_w_data_3 (.hex(reg_w_data[15:12]), .ascii(str_print[1381]));
  hex_to_ascii inst_reg_w_data_2 (.hex(reg_w_data[11:8]), .ascii(str_print[1382]));
  hex_to_ascii inst_reg_w_data_1 (.hex(reg_w_data[7:4]), .ascii(str_print[1383]));
  hex_to_ascii inst_reg_w_data_0 (.hex(reg_w_data[3:0]), .ascii(str_print[1384]));


endmodule //string_to_print
module hex_to_ascii (
  input [3:0] hex,
  output[7:0] ascii
);
  assign ascii = (hex > 4'h9) ? {4'h0, hex} + 8'h37 : {4'h0, hex} + 8'h30;
endmodule
